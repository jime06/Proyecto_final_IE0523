`include "dut1.v"
`include "tester_dut1.v"

module testbench_dut1;

endmodule